**********************************
**** OR2 netlist *****
**********************************
.title OR2

vA A vss pwl(0 0 1n 0 1.01n 0 2n 0 2.01n 1 3n 1 3.01n 1 4n 1)
vB B vss pwl(0 0 1n 0 1.01n 1 2n 1 2.01n 0 3n 0 3.01n 1 4n 1)


** CIRCUIT **


** END CIRCUIT **

.end
