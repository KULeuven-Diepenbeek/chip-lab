**********************************
**** SIMPLE INVERTER netlist *****
**********************************
.title Simple Inverter


** CIRCUIT **

XInv input output vdd vss INVERTER param: multfac='1'

** END CIRCUIT **


.end
